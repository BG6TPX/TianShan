module Top(
  input   clock,
  input   reset
);
endmodule
